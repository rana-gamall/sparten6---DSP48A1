module DSP48A1(A,B,C,D,CARRYIN,M,P,CARRYOUT,CARRYOUTF,CLK,OPMODE,CEA,CEB,CEC,CECARRYIN,CED,CEM,CEOPMODE,CEP
,RSTA,RSTB,RSTC,RSTCARRYIN,RSTD,RSTM,RSTOPMODE,RSTP,BCOUT,PCIN,PCOUT,BCIN);
parameter A0REG  = 1'b0;
parameter A1REG  = 1'b1;
parameter B0REG  = 1'b0;
parameter B1REG  = 1'b1;
parameter CREG   = 1'b1;
parameter DREG   = 1'b1;
parameter MREG   = 1'b1;
parameter PREG   = 1'b1;
parameter OPMODEREG  = 1;
parameter CARRYINREG = 1;
parameter CARRYOUTREG =1;
parameter CARRYINSEL ="OPMODE5";   // "OPMODE5" or "CARRYIN"
parameter B_INPUT   = "DIRECT";    // "DIRECT" or "CASCADE"
parameter RSTTYPE   = "SYNC";      //"SYNC"  or "ASYNC"
input [17:0] A,B,D,BCIN;
input [47:0] PCIN;
input [47:0] C;
input [7:0]OPMODE;
input CARRYIN,CLK,CEA,CEB,CEC,CECARRYIN,CED,CEM,CEOPMODE,CEP;
input RSTA,RSTB,RSTC,RSTCARRYIN,RSTD,RSTM,RSTOPMODE,RSTP;
output [17:0] BCOUT;
output [35:0] M;
output [47:0]PCOUT,P;
output CARRYOUT,CARRYOUTF;
wire [17:0] OUT_B, B0_FINAL,A0_FINAL,D_FINAL,A1_FINAL,OUT_PRE,B1_FINAL,PRE_MUX_RESULT;
wire [47:0] C_FINAL,X_MUX_IN2;
wire [47:0] X_MUX_OUT,Z_MUX_OUT,OUT_POST;
wire [7:0] OPMODE_FINAL;
wire[35:0] multi_result,M_FINAL;
wire CARRY_CASCADE,CARRYIN_FINAL,COUT_POST;
assign BCOUT=B1_FINAL;
assign M=M_FINAL;
assign X_MUX_IN2 ={D_FINAL[11:0] ,A1_FINAL,B1_FINAL};
assign PCOUT=P;
assign CARRYOUTF=CARRYOUT;
reg_MUX #(.N(8),.RSTTYPE(RSTTYPE)) opmode_reg (OPMODE,OPMODEREG,OPMODE_FINAL,CLK,RSTOPMODE,CEOPMODE);
assign OUT_B=(B_INPUT=="DIRECT")? B:
             (B_INPUT=="CASCADE") ? BCIN:0;
reg_MUX #(.N(18),.RSTTYPE(RSTTYPE)) B0_reg (OUT_B,B0REG,B0_FINAL,CLK,RSTB,CEB);
reg_MUX #(.N(18),.RSTTYPE(RSTTYPE)) A0_reg (A,A0REG,A0_FINAL,CLK,RSTA,CEA);
reg_MUX #(.N(18),.RSTTYPE(RSTTYPE)) D0_reg (D,DREG,D_FINAL,CLK,RSTD,CED);
reg_MUX #(.N(48),.RSTTYPE(RSTTYPE)) C0_REG (C,CREG,C_FINAL,CLK,RSTC,CEC);
reg_MUX #(.N(18),.RSTTYPE(RSTTYPE)) A1_reg (A0_FINAL,A1REG,A1_FINAL,CLK,RSTA,CEA);
assign OUT_PRE =(OPMODE_FINAL[6]) ? D_FINAL - B0_FINAL : D_FINAL + B0_FINAL;
assign PRE_MUX_RESULT=(OPMODE_FINAL[4]) ? OUT_PRE :B0_FINAL;
reg_MUX #(.N(18),.RSTTYPE(RSTTYPE)) B1_reg (PRE_MUX_RESULT,B1REG,B1_FINAL,CLK,RSTB,CEB);
assign multi_result =A1_FINAL*B1_FINAL;
reg_MUX #(.N(36),.RSTTYPE(RSTTYPE)) M_reg (multi_result,MREG,M_FINAL,CLK,RSTM,CEM);
MUX4_1 #(.N(48)) X_MUX ({12'h0000,M_FINAL},PCOUT,X_MUX_IN2,OPMODE_FINAL[1:0],X_MUX_OUT);
MUX4_1 #(.N(48)) Z_MUX (PCIN,PCOUT,C_FINAL,OPMODE_FINAL[3:2],Z_MUX_OUT);
assign CARRY_CASCADE =(CARRYINSEL=="OPMODE5") ? OPMODE_FINAL[5]:
                      (CARRYINSEL=="CARRYIN") ? CARRYIN:0;
reg_MUX #(.N(1),.RSTTYPE(RSTTYPE)) carryin_reg (CARRY_CASCADE,CARRYINREG,CARRYIN_FINAL,CLK,RSTCARRYIN,CECARRYIN);
assign {COUT_POST,OUT_POST} =(OPMODE_FINAL[7]) ? Z_MUX_OUT - (X_MUX_OUT + CARRYIN_FINAL) :  Z_MUX_OUT + X_MUX_OUT + CARRYIN_FINAL;
reg_MUX #(.N(48),.RSTTYPE(RSTTYPE)) P_reg (OUT_POST,PREG,P,CLK,RSTP,CEP);
reg_MUX #(.N(1),.RSTTYPE(RSTTYPE)) carryout (COUT_POST,CARRYOUTREG,CARRYOUT,CLK,RSTCARRYIN,CECARRYIN);
endmodule

